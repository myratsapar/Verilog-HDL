modulet lightled(SW, LEDR);
input [17:0] SW;
output [17:0] LEDR;
assign LEDR = SW;
endmodule //3:20 PM 30-Mar-18