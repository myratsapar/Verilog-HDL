module sevenb(HEX0); //b
output [6:0] HEX0;

assign HEX0[0] = 1;
assign HEX0[1] = 1;
assign HEX0[2] = 0;
assign HEX0[3] = 0;
assign HEX0[4] = 0;
assign HEX0[5] = 0;
assign HEX0[6] = 0;

endmodule//7:33 PM 30-Mar-18

